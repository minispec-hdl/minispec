shadowing.ms