lexer1.ms