function4.ms