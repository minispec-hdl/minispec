ctx.ms