function3.ms