function2.ms