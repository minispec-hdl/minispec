function1.ms