function5.ms