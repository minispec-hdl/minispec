lexer2.ms