function Bit#(2) foo(Bit#(2) a, Bit#(2) b) = {a, b};
